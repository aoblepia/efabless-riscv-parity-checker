magic
tech gf180mcuD
magscale 1 5
timestamp 1702248820
<< obsm1 >>
rect 2172 3038 280828 175578
<< metal2 >>
rect 5516 297780 5628 298500
rect 16548 297780 16660 298500
rect 27580 297780 27692 298500
rect 38612 297780 38724 298500
rect 49644 297780 49756 298500
rect 60676 297780 60788 298500
rect 71708 297780 71820 298500
rect 82740 297780 82852 298500
rect 93772 297780 93884 298500
rect 104804 297780 104916 298500
rect 115836 297780 115948 298500
rect 126868 297780 126980 298500
rect 137900 297780 138012 298500
rect 148932 297780 149044 298500
rect 159964 297780 160076 298500
rect 170996 297780 171108 298500
rect 182028 297780 182140 298500
rect 193060 297780 193172 298500
rect 204092 297780 204204 298500
rect 215124 297780 215236 298500
rect 226156 297780 226268 298500
rect 237188 297780 237300 298500
rect 248220 297780 248332 298500
rect 259252 297780 259364 298500
rect 270284 297780 270396 298500
rect 281316 297780 281428 298500
rect 292348 297780 292460 298500
rect 5684 -480 5796 240
rect 6636 -480 6748 240
rect 7588 -480 7700 240
rect 8540 -480 8652 240
rect 9492 -480 9604 240
rect 10444 -480 10556 240
rect 11396 -480 11508 240
rect 12348 -480 12460 240
rect 13300 -480 13412 240
rect 14252 -480 14364 240
rect 15204 -480 15316 240
rect 16156 -480 16268 240
rect 17108 -480 17220 240
rect 18060 -480 18172 240
rect 19012 -480 19124 240
rect 19964 -480 20076 240
rect 20916 -480 21028 240
rect 21868 -480 21980 240
rect 22820 -480 22932 240
rect 23772 -480 23884 240
rect 24724 -480 24836 240
rect 25676 -480 25788 240
rect 26628 -480 26740 240
rect 27580 -480 27692 240
rect 28532 -480 28644 240
rect 29484 -480 29596 240
rect 30436 -480 30548 240
rect 31388 -480 31500 240
rect 32340 -480 32452 240
rect 33292 -480 33404 240
rect 34244 -480 34356 240
rect 35196 -480 35308 240
rect 36148 -480 36260 240
rect 37100 -480 37212 240
rect 38052 -480 38164 240
rect 39004 -480 39116 240
rect 39956 -480 40068 240
rect 40908 -480 41020 240
rect 41860 -480 41972 240
rect 42812 -480 42924 240
rect 43764 -480 43876 240
rect 44716 -480 44828 240
rect 45668 -480 45780 240
rect 46620 -480 46732 240
rect 47572 -480 47684 240
rect 48524 -480 48636 240
rect 49476 -480 49588 240
rect 50428 -480 50540 240
rect 51380 -480 51492 240
rect 52332 -480 52444 240
rect 53284 -480 53396 240
rect 54236 -480 54348 240
rect 55188 -480 55300 240
rect 56140 -480 56252 240
rect 57092 -480 57204 240
rect 58044 -480 58156 240
rect 58996 -480 59108 240
rect 59948 -480 60060 240
rect 60900 -480 61012 240
rect 61852 -480 61964 240
rect 62804 -480 62916 240
rect 63756 -480 63868 240
rect 64708 -480 64820 240
rect 65660 -480 65772 240
rect 66612 -480 66724 240
rect 67564 -480 67676 240
rect 68516 -480 68628 240
rect 69468 -480 69580 240
rect 70420 -480 70532 240
rect 71372 -480 71484 240
rect 72324 -480 72436 240
rect 73276 -480 73388 240
rect 74228 -480 74340 240
rect 75180 -480 75292 240
rect 76132 -480 76244 240
rect 77084 -480 77196 240
rect 78036 -480 78148 240
rect 78988 -480 79100 240
rect 79940 -480 80052 240
rect 80892 -480 81004 240
rect 81844 -480 81956 240
rect 82796 -480 82908 240
rect 83748 -480 83860 240
rect 84700 -480 84812 240
rect 85652 -480 85764 240
rect 86604 -480 86716 240
rect 87556 -480 87668 240
rect 88508 -480 88620 240
rect 89460 -480 89572 240
rect 90412 -480 90524 240
rect 91364 -480 91476 240
rect 92316 -480 92428 240
rect 93268 -480 93380 240
rect 94220 -480 94332 240
rect 95172 -480 95284 240
rect 96124 -480 96236 240
rect 97076 -480 97188 240
rect 98028 -480 98140 240
rect 98980 -480 99092 240
rect 99932 -480 100044 240
rect 100884 -480 100996 240
rect 101836 -480 101948 240
rect 102788 -480 102900 240
rect 103740 -480 103852 240
rect 104692 -480 104804 240
rect 105644 -480 105756 240
rect 106596 -480 106708 240
rect 107548 -480 107660 240
rect 108500 -480 108612 240
rect 109452 -480 109564 240
rect 110404 -480 110516 240
rect 111356 -480 111468 240
rect 112308 -480 112420 240
rect 113260 -480 113372 240
rect 114212 -480 114324 240
rect 115164 -480 115276 240
rect 116116 -480 116228 240
rect 117068 -480 117180 240
rect 118020 -480 118132 240
rect 118972 -480 119084 240
rect 119924 -480 120036 240
rect 120876 -480 120988 240
rect 121828 -480 121940 240
rect 122780 -480 122892 240
rect 123732 -480 123844 240
rect 124684 -480 124796 240
rect 125636 -480 125748 240
rect 126588 -480 126700 240
rect 127540 -480 127652 240
rect 128492 -480 128604 240
rect 129444 -480 129556 240
rect 130396 -480 130508 240
rect 131348 -480 131460 240
rect 132300 -480 132412 240
rect 133252 -480 133364 240
rect 134204 -480 134316 240
rect 135156 -480 135268 240
rect 136108 -480 136220 240
rect 137060 -480 137172 240
rect 138012 -480 138124 240
rect 138964 -480 139076 240
rect 139916 -480 140028 240
rect 140868 -480 140980 240
rect 141820 -480 141932 240
rect 142772 -480 142884 240
rect 143724 -480 143836 240
rect 144676 -480 144788 240
rect 145628 -480 145740 240
rect 146580 -480 146692 240
rect 147532 -480 147644 240
rect 148484 -480 148596 240
rect 149436 -480 149548 240
rect 150388 -480 150500 240
rect 151340 -480 151452 240
rect 152292 -480 152404 240
rect 153244 -480 153356 240
rect 154196 -480 154308 240
rect 155148 -480 155260 240
rect 156100 -480 156212 240
rect 157052 -480 157164 240
rect 158004 -480 158116 240
rect 158956 -480 159068 240
rect 159908 -480 160020 240
rect 160860 -480 160972 240
rect 161812 -480 161924 240
rect 162764 -480 162876 240
rect 163716 -480 163828 240
rect 164668 -480 164780 240
rect 165620 -480 165732 240
rect 166572 -480 166684 240
rect 167524 -480 167636 240
rect 168476 -480 168588 240
rect 169428 -480 169540 240
rect 170380 -480 170492 240
rect 171332 -480 171444 240
rect 172284 -480 172396 240
rect 173236 -480 173348 240
rect 174188 -480 174300 240
rect 175140 -480 175252 240
rect 176092 -480 176204 240
rect 177044 -480 177156 240
rect 177996 -480 178108 240
rect 178948 -480 179060 240
rect 179900 -480 180012 240
rect 180852 -480 180964 240
rect 181804 -480 181916 240
rect 182756 -480 182868 240
rect 183708 -480 183820 240
rect 184660 -480 184772 240
rect 185612 -480 185724 240
rect 186564 -480 186676 240
rect 187516 -480 187628 240
rect 188468 -480 188580 240
rect 189420 -480 189532 240
rect 190372 -480 190484 240
rect 191324 -480 191436 240
rect 192276 -480 192388 240
rect 193228 -480 193340 240
rect 194180 -480 194292 240
rect 195132 -480 195244 240
rect 196084 -480 196196 240
rect 197036 -480 197148 240
rect 197988 -480 198100 240
rect 198940 -480 199052 240
rect 199892 -480 200004 240
rect 200844 -480 200956 240
rect 201796 -480 201908 240
rect 202748 -480 202860 240
rect 203700 -480 203812 240
rect 204652 -480 204764 240
rect 205604 -480 205716 240
rect 206556 -480 206668 240
rect 207508 -480 207620 240
rect 208460 -480 208572 240
rect 209412 -480 209524 240
rect 210364 -480 210476 240
rect 211316 -480 211428 240
rect 212268 -480 212380 240
rect 213220 -480 213332 240
rect 214172 -480 214284 240
rect 215124 -480 215236 240
rect 216076 -480 216188 240
rect 217028 -480 217140 240
rect 217980 -480 218092 240
rect 218932 -480 219044 240
rect 219884 -480 219996 240
rect 220836 -480 220948 240
rect 221788 -480 221900 240
rect 222740 -480 222852 240
rect 223692 -480 223804 240
rect 224644 -480 224756 240
rect 225596 -480 225708 240
rect 226548 -480 226660 240
rect 227500 -480 227612 240
rect 228452 -480 228564 240
rect 229404 -480 229516 240
rect 230356 -480 230468 240
rect 231308 -480 231420 240
rect 232260 -480 232372 240
rect 233212 -480 233324 240
rect 234164 -480 234276 240
rect 235116 -480 235228 240
rect 236068 -480 236180 240
rect 237020 -480 237132 240
rect 237972 -480 238084 240
rect 238924 -480 239036 240
rect 239876 -480 239988 240
rect 240828 -480 240940 240
rect 241780 -480 241892 240
rect 242732 -480 242844 240
rect 243684 -480 243796 240
rect 244636 -480 244748 240
rect 245588 -480 245700 240
rect 246540 -480 246652 240
rect 247492 -480 247604 240
rect 248444 -480 248556 240
rect 249396 -480 249508 240
rect 250348 -480 250460 240
rect 251300 -480 251412 240
rect 252252 -480 252364 240
rect 253204 -480 253316 240
rect 254156 -480 254268 240
rect 255108 -480 255220 240
rect 256060 -480 256172 240
rect 257012 -480 257124 240
rect 257964 -480 258076 240
rect 258916 -480 259028 240
rect 259868 -480 259980 240
rect 260820 -480 260932 240
rect 261772 -480 261884 240
rect 262724 -480 262836 240
rect 263676 -480 263788 240
rect 264628 -480 264740 240
rect 265580 -480 265692 240
rect 266532 -480 266644 240
rect 267484 -480 267596 240
rect 268436 -480 268548 240
rect 269388 -480 269500 240
rect 270340 -480 270452 240
rect 271292 -480 271404 240
rect 272244 -480 272356 240
rect 273196 -480 273308 240
rect 274148 -480 274260 240
rect 275100 -480 275212 240
rect 276052 -480 276164 240
rect 277004 -480 277116 240
rect 277956 -480 278068 240
rect 278908 -480 279020 240
rect 279860 -480 279972 240
rect 280812 -480 280924 240
rect 281764 -480 281876 240
rect 282716 -480 282828 240
rect 283668 -480 283780 240
rect 284620 -480 284732 240
rect 285572 -480 285684 240
rect 286524 -480 286636 240
rect 287476 -480 287588 240
rect 288428 -480 288540 240
rect 289380 -480 289492 240
rect 290332 -480 290444 240
rect 291284 -480 291396 240
rect 292236 -480 292348 240
<< obsm2 >>
rect 2354 297750 5486 297836
rect 5658 297750 16518 297836
rect 16690 297750 27550 297836
rect 27722 297750 38582 297836
rect 38754 297750 49614 297836
rect 49786 297750 60646 297836
rect 60818 297750 71678 297836
rect 71850 297750 82710 297836
rect 82882 297750 93742 297836
rect 93914 297750 104774 297836
rect 104946 297750 115806 297836
rect 115978 297750 126838 297836
rect 127010 297750 137870 297836
rect 138042 297750 148902 297836
rect 149074 297750 159934 297836
rect 160106 297750 170966 297836
rect 171138 297750 181998 297836
rect 182170 297750 193030 297836
rect 193202 297750 204062 297836
rect 204234 297750 215094 297836
rect 215266 297750 226126 297836
rect 226298 297750 237158 297836
rect 237330 297750 248190 297836
rect 248362 297750 259222 297836
rect 259394 297750 270254 297836
rect 270426 297750 281286 297836
rect 281458 297750 282282 297836
rect 2354 270 282282 297750
rect 2354 9 5654 270
rect 5826 9 6606 270
rect 6778 9 7558 270
rect 7730 9 8510 270
rect 8682 9 9462 270
rect 9634 9 10414 270
rect 10586 9 11366 270
rect 11538 9 12318 270
rect 12490 9 13270 270
rect 13442 9 14222 270
rect 14394 9 15174 270
rect 15346 9 16126 270
rect 16298 9 17078 270
rect 17250 9 18030 270
rect 18202 9 18982 270
rect 19154 9 19934 270
rect 20106 9 20886 270
rect 21058 9 21838 270
rect 22010 9 22790 270
rect 22962 9 23742 270
rect 23914 9 24694 270
rect 24866 9 25646 270
rect 25818 9 26598 270
rect 26770 9 27550 270
rect 27722 9 28502 270
rect 28674 9 29454 270
rect 29626 9 30406 270
rect 30578 9 31358 270
rect 31530 9 32310 270
rect 32482 9 33262 270
rect 33434 9 34214 270
rect 34386 9 35166 270
rect 35338 9 36118 270
rect 36290 9 37070 270
rect 37242 9 38022 270
rect 38194 9 38974 270
rect 39146 9 39926 270
rect 40098 9 40878 270
rect 41050 9 41830 270
rect 42002 9 42782 270
rect 42954 9 43734 270
rect 43906 9 44686 270
rect 44858 9 45638 270
rect 45810 9 46590 270
rect 46762 9 47542 270
rect 47714 9 48494 270
rect 48666 9 49446 270
rect 49618 9 50398 270
rect 50570 9 51350 270
rect 51522 9 52302 270
rect 52474 9 53254 270
rect 53426 9 54206 270
rect 54378 9 55158 270
rect 55330 9 56110 270
rect 56282 9 57062 270
rect 57234 9 58014 270
rect 58186 9 58966 270
rect 59138 9 59918 270
rect 60090 9 60870 270
rect 61042 9 61822 270
rect 61994 9 62774 270
rect 62946 9 63726 270
rect 63898 9 64678 270
rect 64850 9 65630 270
rect 65802 9 66582 270
rect 66754 9 67534 270
rect 67706 9 68486 270
rect 68658 9 69438 270
rect 69610 9 70390 270
rect 70562 9 71342 270
rect 71514 9 72294 270
rect 72466 9 73246 270
rect 73418 9 74198 270
rect 74370 9 75150 270
rect 75322 9 76102 270
rect 76274 9 77054 270
rect 77226 9 78006 270
rect 78178 9 78958 270
rect 79130 9 79910 270
rect 80082 9 80862 270
rect 81034 9 81814 270
rect 81986 9 82766 270
rect 82938 9 83718 270
rect 83890 9 84670 270
rect 84842 9 85622 270
rect 85794 9 86574 270
rect 86746 9 87526 270
rect 87698 9 88478 270
rect 88650 9 89430 270
rect 89602 9 90382 270
rect 90554 9 91334 270
rect 91506 9 92286 270
rect 92458 9 93238 270
rect 93410 9 94190 270
rect 94362 9 95142 270
rect 95314 9 96094 270
rect 96266 9 97046 270
rect 97218 9 97998 270
rect 98170 9 98950 270
rect 99122 9 99902 270
rect 100074 9 100854 270
rect 101026 9 101806 270
rect 101978 9 102758 270
rect 102930 9 103710 270
rect 103882 9 104662 270
rect 104834 9 105614 270
rect 105786 9 106566 270
rect 106738 9 107518 270
rect 107690 9 108470 270
rect 108642 9 109422 270
rect 109594 9 110374 270
rect 110546 9 111326 270
rect 111498 9 112278 270
rect 112450 9 113230 270
rect 113402 9 114182 270
rect 114354 9 115134 270
rect 115306 9 116086 270
rect 116258 9 117038 270
rect 117210 9 117990 270
rect 118162 9 118942 270
rect 119114 9 119894 270
rect 120066 9 120846 270
rect 121018 9 121798 270
rect 121970 9 122750 270
rect 122922 9 123702 270
rect 123874 9 124654 270
rect 124826 9 125606 270
rect 125778 9 126558 270
rect 126730 9 127510 270
rect 127682 9 128462 270
rect 128634 9 129414 270
rect 129586 9 130366 270
rect 130538 9 131318 270
rect 131490 9 132270 270
rect 132442 9 133222 270
rect 133394 9 134174 270
rect 134346 9 135126 270
rect 135298 9 136078 270
rect 136250 9 137030 270
rect 137202 9 137982 270
rect 138154 9 138934 270
rect 139106 9 139886 270
rect 140058 9 140838 270
rect 141010 9 141790 270
rect 141962 9 142742 270
rect 142914 9 143694 270
rect 143866 9 144646 270
rect 144818 9 145598 270
rect 145770 9 146550 270
rect 146722 9 147502 270
rect 147674 9 148454 270
rect 148626 9 149406 270
rect 149578 9 150358 270
rect 150530 9 151310 270
rect 151482 9 152262 270
rect 152434 9 153214 270
rect 153386 9 154166 270
rect 154338 9 155118 270
rect 155290 9 156070 270
rect 156242 9 157022 270
rect 157194 9 157974 270
rect 158146 9 158926 270
rect 159098 9 159878 270
rect 160050 9 160830 270
rect 161002 9 161782 270
rect 161954 9 162734 270
rect 162906 9 163686 270
rect 163858 9 164638 270
rect 164810 9 165590 270
rect 165762 9 166542 270
rect 166714 9 167494 270
rect 167666 9 168446 270
rect 168618 9 169398 270
rect 169570 9 170350 270
rect 170522 9 171302 270
rect 171474 9 172254 270
rect 172426 9 173206 270
rect 173378 9 174158 270
rect 174330 9 175110 270
rect 175282 9 176062 270
rect 176234 9 177014 270
rect 177186 9 177966 270
rect 178138 9 178918 270
rect 179090 9 179870 270
rect 180042 9 180822 270
rect 180994 9 181774 270
rect 181946 9 182726 270
rect 182898 9 183678 270
rect 183850 9 184630 270
rect 184802 9 185582 270
rect 185754 9 186534 270
rect 186706 9 187486 270
rect 187658 9 188438 270
rect 188610 9 189390 270
rect 189562 9 190342 270
rect 190514 9 191294 270
rect 191466 9 192246 270
rect 192418 9 193198 270
rect 193370 9 194150 270
rect 194322 9 195102 270
rect 195274 9 196054 270
rect 196226 9 197006 270
rect 197178 9 197958 270
rect 198130 9 198910 270
rect 199082 9 199862 270
rect 200034 9 200814 270
rect 200986 9 201766 270
rect 201938 9 202718 270
rect 202890 9 203670 270
rect 203842 9 204622 270
rect 204794 9 205574 270
rect 205746 9 206526 270
rect 206698 9 207478 270
rect 207650 9 208430 270
rect 208602 9 209382 270
rect 209554 9 210334 270
rect 210506 9 211286 270
rect 211458 9 212238 270
rect 212410 9 213190 270
rect 213362 9 214142 270
rect 214314 9 215094 270
rect 215266 9 216046 270
rect 216218 9 216998 270
rect 217170 9 217950 270
rect 218122 9 218902 270
rect 219074 9 219854 270
rect 220026 9 220806 270
rect 220978 9 221758 270
rect 221930 9 222710 270
rect 222882 9 223662 270
rect 223834 9 224614 270
rect 224786 9 225566 270
rect 225738 9 226518 270
rect 226690 9 227470 270
rect 227642 9 228422 270
rect 228594 9 229374 270
rect 229546 9 230326 270
rect 230498 9 231278 270
rect 231450 9 232230 270
rect 232402 9 233182 270
rect 233354 9 234134 270
rect 234306 9 235086 270
rect 235258 9 236038 270
rect 236210 9 236990 270
rect 237162 9 237942 270
rect 238114 9 238894 270
rect 239066 9 239846 270
rect 240018 9 240798 270
rect 240970 9 241750 270
rect 241922 9 242702 270
rect 242874 9 243654 270
rect 243826 9 244606 270
rect 244778 9 245558 270
rect 245730 9 246510 270
rect 246682 9 247462 270
rect 247634 9 248414 270
rect 248586 9 249366 270
rect 249538 9 250318 270
rect 250490 9 251270 270
rect 251442 9 252222 270
rect 252394 9 253174 270
rect 253346 9 254126 270
rect 254298 9 255078 270
rect 255250 9 256030 270
rect 256202 9 256982 270
rect 257154 9 257934 270
rect 258106 9 258886 270
rect 259058 9 259838 270
rect 260010 9 260790 270
rect 260962 9 261742 270
rect 261914 9 262694 270
rect 262866 9 263646 270
rect 263818 9 264598 270
rect 264770 9 265550 270
rect 265722 9 266502 270
rect 266674 9 267454 270
rect 267626 9 268406 270
rect 268578 9 269358 270
rect 269530 9 270310 270
rect 270482 9 271262 270
rect 271434 9 272214 270
rect 272386 9 273166 270
rect 273338 9 274118 270
rect 274290 9 275070 270
rect 275242 9 276022 270
rect 276194 9 276974 270
rect 277146 9 277926 270
rect 278098 9 278878 270
rect 279050 9 279830 270
rect 280002 9 280782 270
rect 280954 9 281734 270
rect 281906 9 282282 270
<< metal3 >>
rect 297780 294308 298500 294420
rect -480 293580 240 293692
rect 297780 287700 298500 287812
rect -480 286524 240 286636
rect 297780 281092 298500 281204
rect -480 279468 240 279580
rect 297780 274484 298500 274596
rect -480 272412 240 272524
rect 297780 267876 298500 267988
rect -480 265356 240 265468
rect 297780 261268 298500 261380
rect -480 258300 240 258412
rect 297780 254660 298500 254772
rect -480 251244 240 251356
rect 297780 248052 298500 248164
rect -480 244188 240 244300
rect 297780 241444 298500 241556
rect -480 237132 240 237244
rect 297780 234836 298500 234948
rect -480 230076 240 230188
rect 297780 228228 298500 228340
rect -480 223020 240 223132
rect 297780 221620 298500 221732
rect -480 215964 240 216076
rect 297780 215012 298500 215124
rect -480 208908 240 209020
rect 297780 208404 298500 208516
rect -480 201852 240 201964
rect 297780 201796 298500 201908
rect 297780 195188 298500 195300
rect -480 194796 240 194908
rect 297780 188580 298500 188692
rect -480 187740 240 187852
rect 297780 181972 298500 182084
rect -480 180684 240 180796
rect 297780 175364 298500 175476
rect -480 173628 240 173740
rect 297780 168756 298500 168868
rect -480 166572 240 166684
rect 297780 162148 298500 162260
rect -480 159516 240 159628
rect 297780 155540 298500 155652
rect -480 152460 240 152572
rect 297780 148932 298500 149044
rect -480 145404 240 145516
rect 297780 142324 298500 142436
rect -480 138348 240 138460
rect 297780 135716 298500 135828
rect -480 131292 240 131404
rect 297780 129108 298500 129220
rect -480 124236 240 124348
rect 297780 122500 298500 122612
rect -480 117180 240 117292
rect 297780 115892 298500 116004
rect -480 110124 240 110236
rect 297780 109284 298500 109396
rect -480 103068 240 103180
rect 297780 102676 298500 102788
rect -480 96012 240 96124
rect 297780 96068 298500 96180
rect 297780 89460 298500 89572
rect -480 88956 240 89068
rect 297780 82852 298500 82964
rect -480 81900 240 82012
rect 297780 76244 298500 76356
rect -480 74844 240 74956
rect 297780 69636 298500 69748
rect -480 67788 240 67900
rect 297780 63028 298500 63140
rect -480 60732 240 60844
rect 297780 56420 298500 56532
rect -480 53676 240 53788
rect 297780 49812 298500 49924
rect -480 46620 240 46732
rect 297780 43204 298500 43316
rect -480 39564 240 39676
rect 297780 36596 298500 36708
rect -480 32508 240 32620
rect 297780 29988 298500 30100
rect -480 25452 240 25564
rect 297780 23380 298500 23492
rect -480 18396 240 18508
rect 297780 16772 298500 16884
rect -480 11340 240 11452
rect 297780 10164 298500 10276
rect -480 4284 240 4396
rect 297780 3556 298500 3668
<< obsm3 >>
rect 793 294450 297836 295330
rect 793 294278 297750 294450
rect 793 287842 297836 294278
rect 793 287670 297750 287842
rect 793 281234 297836 287670
rect 793 281062 297750 281234
rect 793 274626 297836 281062
rect 793 274454 297750 274626
rect 793 268018 297836 274454
rect 793 267846 297750 268018
rect 793 261410 297836 267846
rect 793 261238 297750 261410
rect 793 254802 297836 261238
rect 793 254630 297750 254802
rect 793 248194 297836 254630
rect 793 248022 297750 248194
rect 793 241586 297836 248022
rect 793 241414 297750 241586
rect 793 234978 297836 241414
rect 793 234806 297750 234978
rect 793 228370 297836 234806
rect 793 228198 297750 228370
rect 793 221762 297836 228198
rect 793 221590 297750 221762
rect 793 215154 297836 221590
rect 793 214982 297750 215154
rect 793 208546 297836 214982
rect 793 208374 297750 208546
rect 793 201938 297836 208374
rect 793 201766 297750 201938
rect 793 195330 297836 201766
rect 793 195158 297750 195330
rect 793 188722 297836 195158
rect 793 188550 297750 188722
rect 793 182114 297836 188550
rect 793 181942 297750 182114
rect 793 175506 297836 181942
rect 793 175334 297750 175506
rect 793 168898 297836 175334
rect 793 168726 297750 168898
rect 793 162290 297836 168726
rect 793 162118 297750 162290
rect 793 155682 297836 162118
rect 793 155510 297750 155682
rect 793 149074 297836 155510
rect 793 148902 297750 149074
rect 793 142466 297836 148902
rect 793 142294 297750 142466
rect 793 135858 297836 142294
rect 793 135686 297750 135858
rect 793 129250 297836 135686
rect 793 129078 297750 129250
rect 793 122642 297836 129078
rect 793 122470 297750 122642
rect 793 116034 297836 122470
rect 793 115862 297750 116034
rect 793 109426 297836 115862
rect 793 109254 297750 109426
rect 793 102818 297836 109254
rect 793 102646 297750 102818
rect 793 96210 297836 102646
rect 793 96038 297750 96210
rect 793 89602 297836 96038
rect 793 89430 297750 89602
rect 793 82994 297836 89430
rect 793 82822 297750 82994
rect 793 76386 297836 82822
rect 793 76214 297750 76386
rect 793 69778 297836 76214
rect 793 69606 297750 69778
rect 793 63170 297836 69606
rect 793 62998 297750 63170
rect 793 56562 297836 62998
rect 793 56390 297750 56562
rect 793 49954 297836 56390
rect 793 49782 297750 49954
rect 793 43346 297836 49782
rect 793 43174 297750 43346
rect 793 36738 297836 43174
rect 793 36566 297750 36738
rect 793 30130 297836 36566
rect 793 29958 297750 30130
rect 793 23522 297836 29958
rect 793 23350 297750 23522
rect 793 16914 297836 23350
rect 793 16742 297750 16914
rect 793 10306 297836 16742
rect 793 10134 297750 10306
rect 793 3698 297836 10134
rect 793 3526 297750 3698
rect 793 14 297836 3526
<< metal4 >>
rect -958 -822 -648 299134
rect -478 -342 -168 298654
rect 2709 -822 3019 299134
rect 4569 -822 4879 299134
rect 18069 -822 18379 299134
rect 19929 -822 20239 299134
rect 33429 -822 33739 299134
rect 35289 -822 35599 299134
rect 48789 -822 49099 299134
rect 50649 -822 50959 299134
rect 64149 -822 64459 299134
rect 66009 -822 66319 299134
rect 79509 -822 79819 299134
rect 81369 -822 81679 299134
rect 94869 -822 95179 299134
rect 96729 -822 97039 299134
rect 110229 -822 110539 299134
rect 112089 -822 112399 299134
rect 125589 -822 125899 299134
rect 127449 -822 127759 299134
rect 140949 -822 141259 299134
rect 142809 -822 143119 299134
rect 156309 -822 156619 299134
rect 158169 -822 158479 299134
rect 171669 -822 171979 299134
rect 173529 -822 173839 299134
rect 187029 -822 187339 299134
rect 188889 -822 189199 299134
rect 202389 -822 202699 299134
rect 204249 -822 204559 299134
rect 217749 -822 218059 299134
rect 219609 -822 219919 299134
rect 233109 -822 233419 299134
rect 234969 -822 235279 299134
rect 248469 -822 248779 299134
rect 250329 -822 250639 299134
rect 263829 -822 264139 299134
rect 265689 -822 265999 299134
rect 279189 -822 279499 299134
rect 281049 112587 281359 299134
rect 281049 -822 281359 109205
rect 294549 -822 294859 299134
rect 296409 -822 296719 299134
rect 298200 -342 298510 298654
rect 298680 -822 298990 299134
<< obsm4 >>
rect 798 3038 2679 295111
rect 3049 3038 4539 295111
rect 4909 3038 18039 295111
rect 18409 3038 19899 295111
rect 20269 3038 33399 295111
rect 33769 3038 35259 295111
rect 35629 3038 48759 295111
rect 49129 3038 50619 295111
rect 50989 3038 64119 295111
rect 64489 3038 65979 295111
rect 66349 3038 79479 295111
rect 79849 3038 81339 295111
rect 81709 3038 94839 295111
rect 95209 3038 96699 295111
rect 97069 3038 110199 295111
rect 110569 3038 112059 295111
rect 112429 3038 125559 295111
rect 125929 3038 127419 295111
rect 127789 3038 140919 295111
rect 141289 3038 142779 295111
rect 143149 3038 156279 295111
rect 156649 3038 158139 295111
rect 158509 3038 171639 295111
rect 172009 3038 173499 295111
rect 173869 3038 186999 295111
rect 187369 3038 188859 295111
rect 189229 3038 202359 295111
rect 202729 3038 204219 295111
rect 204589 3038 217719 295111
rect 218089 3038 219579 295111
rect 219949 3038 233079 295111
rect 233449 3038 234939 295111
rect 235309 3038 248439 295111
rect 248809 3038 250299 295111
rect 250669 3038 263799 295111
rect 264169 3038 265659 295111
rect 266029 3038 279159 295111
rect 279529 112557 281019 295111
rect 281389 112557 294519 295111
rect 279529 109235 294519 112557
rect 279529 3038 281019 109235
rect 281389 3038 294519 109235
rect 294889 3038 295330 295111
<< metal5 >>
rect -958 298824 298990 299134
rect -478 298344 298510 298654
rect -958 292913 298990 293223
rect -958 289913 298990 290223
rect -958 283913 298990 284223
rect -958 280913 298990 281223
rect -958 274913 298990 275223
rect -958 271913 298990 272223
rect -958 265913 298990 266223
rect -958 262913 298990 263223
rect -958 256913 298990 257223
rect -958 253913 298990 254223
rect -958 247913 298990 248223
rect -958 244913 298990 245223
rect -958 238913 298990 239223
rect -958 235913 298990 236223
rect -958 229913 298990 230223
rect -958 226913 298990 227223
rect -958 220913 298990 221223
rect -958 217913 298990 218223
rect -958 211913 298990 212223
rect -958 208913 298990 209223
rect -958 202913 298990 203223
rect -958 199913 298990 200223
rect -958 193913 298990 194223
rect -958 190913 298990 191223
rect -958 184913 298990 185223
rect -958 181913 298990 182223
rect -958 175913 298990 176223
rect -958 172913 298990 173223
rect -958 166913 298990 167223
rect -958 163913 298990 164223
rect -958 157913 298990 158223
rect -958 154913 298990 155223
rect -958 148913 298990 149223
rect -958 145913 298990 146223
rect -958 139913 298990 140223
rect -958 136913 298990 137223
rect -958 130913 298990 131223
rect -958 127913 298990 128223
rect -958 121913 298990 122223
rect -958 118913 298990 119223
rect -958 112913 298990 113223
rect -958 109913 298990 110223
rect -958 103913 298990 104223
rect -958 100913 298990 101223
rect -958 94913 298990 95223
rect -958 91913 298990 92223
rect -958 85913 298990 86223
rect -958 82913 298990 83223
rect -958 76913 298990 77223
rect -958 73913 298990 74223
rect -958 67913 298990 68223
rect -958 64913 298990 65223
rect -958 58913 298990 59223
rect -958 55913 298990 56223
rect -958 49913 298990 50223
rect -958 46913 298990 47223
rect -958 40913 298990 41223
rect -958 37913 298990 38223
rect -958 31913 298990 32223
rect -958 28913 298990 29223
rect -958 22913 298990 23223
rect -958 19913 298990 20223
rect -958 13913 298990 14223
rect -958 10913 298990 11223
rect -958 4913 298990 5223
rect -958 1913 298990 2223
rect -478 -342 298510 -32
rect -958 -822 298990 -512
<< obsm5 >>
rect 248366 95693 281450 95737
<< labels >>
rlabel metal3 s 297780 3556 298500 3668 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 297780 201796 298500 201908 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 297780 221620 298500 221732 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 297780 241444 298500 241556 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 297780 261268 298500 261380 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 297780 281092 298500 281204 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 292348 297780 292460 298500 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 259252 297780 259364 298500 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 226156 297780 226268 298500 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 193060 297780 193172 298500 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 159964 297780 160076 298500 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 297780 23380 298500 23492 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 126868 297780 126980 298500 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 93772 297780 93884 298500 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 60676 297780 60788 298500 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 27580 297780 27692 298500 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s -480 293580 240 293692 4 io_in[24]
port 17 nsew signal input
rlabel metal3 s -480 272412 240 272524 4 io_in[25]
port 18 nsew signal input
rlabel metal3 s -480 251244 240 251356 4 io_in[26]
port 19 nsew signal input
rlabel metal3 s -480 230076 240 230188 4 io_in[27]
port 20 nsew signal input
rlabel metal3 s -480 208908 240 209020 4 io_in[28]
port 21 nsew signal input
rlabel metal3 s -480 187740 240 187852 4 io_in[29]
port 22 nsew signal input
rlabel metal3 s 297780 43204 298500 43316 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s -480 166572 240 166684 4 io_in[30]
port 24 nsew signal input
rlabel metal3 s -480 145404 240 145516 4 io_in[31]
port 25 nsew signal input
rlabel metal3 s -480 124236 240 124348 4 io_in[32]
port 26 nsew signal input
rlabel metal3 s -480 103068 240 103180 4 io_in[33]
port 27 nsew signal input
rlabel metal3 s -480 81900 240 82012 4 io_in[34]
port 28 nsew signal input
rlabel metal3 s -480 60732 240 60844 4 io_in[35]
port 29 nsew signal input
rlabel metal3 s -480 39564 240 39676 4 io_in[36]
port 30 nsew signal input
rlabel metal3 s -480 18396 240 18508 4 io_in[37]
port 31 nsew signal input
rlabel metal3 s 297780 63028 298500 63140 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 297780 82852 298500 82964 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 297780 102676 298500 102788 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 297780 122500 298500 122612 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 297780 142324 298500 142436 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 297780 162148 298500 162260 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 297780 181972 298500 182084 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 297780 16772 298500 16884 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 297780 215012 298500 215124 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 297780 234836 298500 234948 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 297780 254660 298500 254772 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 297780 274484 298500 274596 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 297780 294308 298500 294420 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 270284 297780 270396 298500 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 237188 297780 237300 298500 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 204092 297780 204204 298500 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 170996 297780 171108 298500 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 137900 297780 138012 298500 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 297780 36596 298500 36708 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 104804 297780 104916 298500 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 71708 297780 71820 298500 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 38612 297780 38724 298500 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 5516 297780 5628 298500 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s -480 279468 240 279580 4 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s -480 258300 240 258412 4 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s -480 237132 240 237244 4 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s -480 215964 240 216076 4 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s -480 194796 240 194908 4 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s -480 173628 240 173740 4 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 297780 56420 298500 56532 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s -480 152460 240 152572 4 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s -480 131292 240 131404 4 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s -480 110124 240 110236 4 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s -480 88956 240 89068 4 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s -480 67788 240 67900 4 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s -480 46620 240 46732 4 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s -480 25452 240 25564 4 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s -480 4284 240 4396 4 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 297780 76244 298500 76356 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 297780 96068 298500 96180 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 297780 115892 298500 116004 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 297780 135716 298500 135828 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 297780 155540 298500 155652 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 297780 175364 298500 175476 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 297780 195188 298500 195300 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 297780 10164 298500 10276 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 297780 208404 298500 208516 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 297780 228228 298500 228340 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 297780 248052 298500 248164 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 297780 267876 298500 267988 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 297780 287700 298500 287812 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 281316 297780 281428 298500 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 248220 297780 248332 298500 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 215124 297780 215236 298500 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 182028 297780 182140 298500 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 148932 297780 149044 298500 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 297780 29988 298500 30100 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 115836 297780 115948 298500 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 82740 297780 82852 298500 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 49644 297780 49756 298500 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 16548 297780 16660 298500 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s -480 286524 240 286636 4 io_out[24]
port 93 nsew signal output
rlabel metal3 s -480 265356 240 265468 4 io_out[25]
port 94 nsew signal output
rlabel metal3 s -480 244188 240 244300 4 io_out[26]
port 95 nsew signal output
rlabel metal3 s -480 223020 240 223132 4 io_out[27]
port 96 nsew signal output
rlabel metal3 s -480 201852 240 201964 4 io_out[28]
port 97 nsew signal output
rlabel metal3 s -480 180684 240 180796 4 io_out[29]
port 98 nsew signal output
rlabel metal3 s 297780 49812 298500 49924 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s -480 159516 240 159628 4 io_out[30]
port 100 nsew signal output
rlabel metal3 s -480 138348 240 138460 4 io_out[31]
port 101 nsew signal output
rlabel metal3 s -480 117180 240 117292 4 io_out[32]
port 102 nsew signal output
rlabel metal3 s -480 96012 240 96124 4 io_out[33]
port 103 nsew signal output
rlabel metal3 s -480 74844 240 74956 4 io_out[34]
port 104 nsew signal output
rlabel metal3 s -480 53676 240 53788 4 io_out[35]
port 105 nsew signal output
rlabel metal3 s -480 32508 240 32620 4 io_out[36]
port 106 nsew signal output
rlabel metal3 s -480 11340 240 11452 4 io_out[37]
port 107 nsew signal output
rlabel metal3 s 297780 69636 298500 69748 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 297780 89460 298500 89572 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 297780 109284 298500 109396 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 297780 129108 298500 129220 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 297780 148932 298500 149044 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 297780 168756 298500 168868 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 297780 188580 298500 188692 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 106596 -480 106708 240 8 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 135156 -480 135268 240 8 la_data_in[10]
port 116 nsew signal input
rlabel metal2 s 138012 -480 138124 240 8 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 140868 -480 140980 240 8 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 143724 -480 143836 240 8 la_data_in[13]
port 119 nsew signal input
rlabel metal2 s 146580 -480 146692 240 8 la_data_in[14]
port 120 nsew signal input
rlabel metal2 s 149436 -480 149548 240 8 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 152292 -480 152404 240 8 la_data_in[16]
port 122 nsew signal input
rlabel metal2 s 155148 -480 155260 240 8 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 158004 -480 158116 240 8 la_data_in[18]
port 124 nsew signal input
rlabel metal2 s 160860 -480 160972 240 8 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 109452 -480 109564 240 8 la_data_in[1]
port 126 nsew signal input
rlabel metal2 s 163716 -480 163828 240 8 la_data_in[20]
port 127 nsew signal input
rlabel metal2 s 166572 -480 166684 240 8 la_data_in[21]
port 128 nsew signal input
rlabel metal2 s 169428 -480 169540 240 8 la_data_in[22]
port 129 nsew signal input
rlabel metal2 s 172284 -480 172396 240 8 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 175140 -480 175252 240 8 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 177996 -480 178108 240 8 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 180852 -480 180964 240 8 la_data_in[26]
port 133 nsew signal input
rlabel metal2 s 183708 -480 183820 240 8 la_data_in[27]
port 134 nsew signal input
rlabel metal2 s 186564 -480 186676 240 8 la_data_in[28]
port 135 nsew signal input
rlabel metal2 s 189420 -480 189532 240 8 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 112308 -480 112420 240 8 la_data_in[2]
port 137 nsew signal input
rlabel metal2 s 192276 -480 192388 240 8 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 195132 -480 195244 240 8 la_data_in[31]
port 139 nsew signal input
rlabel metal2 s 197988 -480 198100 240 8 la_data_in[32]
port 140 nsew signal input
rlabel metal2 s 200844 -480 200956 240 8 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 203700 -480 203812 240 8 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 206556 -480 206668 240 8 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 209412 -480 209524 240 8 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 212268 -480 212380 240 8 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 215124 -480 215236 240 8 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 217980 -480 218092 240 8 la_data_in[39]
port 147 nsew signal input
rlabel metal2 s 115164 -480 115276 240 8 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 220836 -480 220948 240 8 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 223692 -480 223804 240 8 la_data_in[41]
port 150 nsew signal input
rlabel metal2 s 226548 -480 226660 240 8 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 229404 -480 229516 240 8 la_data_in[43]
port 152 nsew signal input
rlabel metal2 s 232260 -480 232372 240 8 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 235116 -480 235228 240 8 la_data_in[45]
port 154 nsew signal input
rlabel metal2 s 237972 -480 238084 240 8 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 240828 -480 240940 240 8 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 243684 -480 243796 240 8 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 246540 -480 246652 240 8 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 118020 -480 118132 240 8 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 249396 -480 249508 240 8 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 252252 -480 252364 240 8 la_data_in[51]
port 161 nsew signal input
rlabel metal2 s 255108 -480 255220 240 8 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 257964 -480 258076 240 8 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 260820 -480 260932 240 8 la_data_in[54]
port 164 nsew signal input
rlabel metal2 s 263676 -480 263788 240 8 la_data_in[55]
port 165 nsew signal input
rlabel metal2 s 266532 -480 266644 240 8 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 269388 -480 269500 240 8 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 272244 -480 272356 240 8 la_data_in[58]
port 168 nsew signal input
rlabel metal2 s 275100 -480 275212 240 8 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 120876 -480 120988 240 8 la_data_in[5]
port 170 nsew signal input
rlabel metal2 s 277956 -480 278068 240 8 la_data_in[60]
port 171 nsew signal input
rlabel metal2 s 280812 -480 280924 240 8 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 283668 -480 283780 240 8 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 286524 -480 286636 240 8 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 123732 -480 123844 240 8 la_data_in[6]
port 175 nsew signal input
rlabel metal2 s 126588 -480 126700 240 8 la_data_in[7]
port 176 nsew signal input
rlabel metal2 s 129444 -480 129556 240 8 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 132300 -480 132412 240 8 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 107548 -480 107660 240 8 la_data_out[0]
port 179 nsew signal output
rlabel metal2 s 136108 -480 136220 240 8 la_data_out[10]
port 180 nsew signal output
rlabel metal2 s 138964 -480 139076 240 8 la_data_out[11]
port 181 nsew signal output
rlabel metal2 s 141820 -480 141932 240 8 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 144676 -480 144788 240 8 la_data_out[13]
port 183 nsew signal output
rlabel metal2 s 147532 -480 147644 240 8 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 150388 -480 150500 240 8 la_data_out[15]
port 185 nsew signal output
rlabel metal2 s 153244 -480 153356 240 8 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 156100 -480 156212 240 8 la_data_out[17]
port 187 nsew signal output
rlabel metal2 s 158956 -480 159068 240 8 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 161812 -480 161924 240 8 la_data_out[19]
port 189 nsew signal output
rlabel metal2 s 110404 -480 110516 240 8 la_data_out[1]
port 190 nsew signal output
rlabel metal2 s 164668 -480 164780 240 8 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 167524 -480 167636 240 8 la_data_out[21]
port 192 nsew signal output
rlabel metal2 s 170380 -480 170492 240 8 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 173236 -480 173348 240 8 la_data_out[23]
port 194 nsew signal output
rlabel metal2 s 176092 -480 176204 240 8 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 178948 -480 179060 240 8 la_data_out[25]
port 196 nsew signal output
rlabel metal2 s 181804 -480 181916 240 8 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 184660 -480 184772 240 8 la_data_out[27]
port 198 nsew signal output
rlabel metal2 s 187516 -480 187628 240 8 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 190372 -480 190484 240 8 la_data_out[29]
port 200 nsew signal output
rlabel metal2 s 113260 -480 113372 240 8 la_data_out[2]
port 201 nsew signal output
rlabel metal2 s 193228 -480 193340 240 8 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 196084 -480 196196 240 8 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 198940 -480 199052 240 8 la_data_out[32]
port 204 nsew signal output
rlabel metal2 s 201796 -480 201908 240 8 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 204652 -480 204764 240 8 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 207508 -480 207620 240 8 la_data_out[35]
port 207 nsew signal output
rlabel metal2 s 210364 -480 210476 240 8 la_data_out[36]
port 208 nsew signal output
rlabel metal2 s 213220 -480 213332 240 8 la_data_out[37]
port 209 nsew signal output
rlabel metal2 s 216076 -480 216188 240 8 la_data_out[38]
port 210 nsew signal output
rlabel metal2 s 218932 -480 219044 240 8 la_data_out[39]
port 211 nsew signal output
rlabel metal2 s 116116 -480 116228 240 8 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 221788 -480 221900 240 8 la_data_out[40]
port 213 nsew signal output
rlabel metal2 s 224644 -480 224756 240 8 la_data_out[41]
port 214 nsew signal output
rlabel metal2 s 227500 -480 227612 240 8 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 230356 -480 230468 240 8 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 233212 -480 233324 240 8 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 236068 -480 236180 240 8 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 238924 -480 239036 240 8 la_data_out[46]
port 219 nsew signal output
rlabel metal2 s 241780 -480 241892 240 8 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 244636 -480 244748 240 8 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 247492 -480 247604 240 8 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 118972 -480 119084 240 8 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 250348 -480 250460 240 8 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 253204 -480 253316 240 8 la_data_out[51]
port 225 nsew signal output
rlabel metal2 s 256060 -480 256172 240 8 la_data_out[52]
port 226 nsew signal output
rlabel metal2 s 258916 -480 259028 240 8 la_data_out[53]
port 227 nsew signal output
rlabel metal2 s 261772 -480 261884 240 8 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 264628 -480 264740 240 8 la_data_out[55]
port 229 nsew signal output
rlabel metal2 s 267484 -480 267596 240 8 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 270340 -480 270452 240 8 la_data_out[57]
port 231 nsew signal output
rlabel metal2 s 273196 -480 273308 240 8 la_data_out[58]
port 232 nsew signal output
rlabel metal2 s 276052 -480 276164 240 8 la_data_out[59]
port 233 nsew signal output
rlabel metal2 s 121828 -480 121940 240 8 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 278908 -480 279020 240 8 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 281764 -480 281876 240 8 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 284620 -480 284732 240 8 la_data_out[62]
port 237 nsew signal output
rlabel metal2 s 287476 -480 287588 240 8 la_data_out[63]
port 238 nsew signal output
rlabel metal2 s 124684 -480 124796 240 8 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 127540 -480 127652 240 8 la_data_out[7]
port 240 nsew signal output
rlabel metal2 s 130396 -480 130508 240 8 la_data_out[8]
port 241 nsew signal output
rlabel metal2 s 133252 -480 133364 240 8 la_data_out[9]
port 242 nsew signal output
rlabel metal2 s 108500 -480 108612 240 8 la_oenb[0]
port 243 nsew signal input
rlabel metal2 s 137060 -480 137172 240 8 la_oenb[10]
port 244 nsew signal input
rlabel metal2 s 139916 -480 140028 240 8 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 142772 -480 142884 240 8 la_oenb[12]
port 246 nsew signal input
rlabel metal2 s 145628 -480 145740 240 8 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 148484 -480 148596 240 8 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 151340 -480 151452 240 8 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 154196 -480 154308 240 8 la_oenb[16]
port 250 nsew signal input
rlabel metal2 s 157052 -480 157164 240 8 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 159908 -480 160020 240 8 la_oenb[18]
port 252 nsew signal input
rlabel metal2 s 162764 -480 162876 240 8 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 111356 -480 111468 240 8 la_oenb[1]
port 254 nsew signal input
rlabel metal2 s 165620 -480 165732 240 8 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 168476 -480 168588 240 8 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 171332 -480 171444 240 8 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 174188 -480 174300 240 8 la_oenb[23]
port 258 nsew signal input
rlabel metal2 s 177044 -480 177156 240 8 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 179900 -480 180012 240 8 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 182756 -480 182868 240 8 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 185612 -480 185724 240 8 la_oenb[27]
port 262 nsew signal input
rlabel metal2 s 188468 -480 188580 240 8 la_oenb[28]
port 263 nsew signal input
rlabel metal2 s 191324 -480 191436 240 8 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 114212 -480 114324 240 8 la_oenb[2]
port 265 nsew signal input
rlabel metal2 s 194180 -480 194292 240 8 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 197036 -480 197148 240 8 la_oenb[31]
port 267 nsew signal input
rlabel metal2 s 199892 -480 200004 240 8 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 202748 -480 202860 240 8 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 205604 -480 205716 240 8 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 208460 -480 208572 240 8 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 211316 -480 211428 240 8 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 214172 -480 214284 240 8 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 217028 -480 217140 240 8 la_oenb[38]
port 274 nsew signal input
rlabel metal2 s 219884 -480 219996 240 8 la_oenb[39]
port 275 nsew signal input
rlabel metal2 s 117068 -480 117180 240 8 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 222740 -480 222852 240 8 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 225596 -480 225708 240 8 la_oenb[41]
port 278 nsew signal input
rlabel metal2 s 228452 -480 228564 240 8 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 231308 -480 231420 240 8 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 234164 -480 234276 240 8 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 237020 -480 237132 240 8 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 239876 -480 239988 240 8 la_oenb[46]
port 283 nsew signal input
rlabel metal2 s 242732 -480 242844 240 8 la_oenb[47]
port 284 nsew signal input
rlabel metal2 s 245588 -480 245700 240 8 la_oenb[48]
port 285 nsew signal input
rlabel metal2 s 248444 -480 248556 240 8 la_oenb[49]
port 286 nsew signal input
rlabel metal2 s 119924 -480 120036 240 8 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 251300 -480 251412 240 8 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 254156 -480 254268 240 8 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 257012 -480 257124 240 8 la_oenb[52]
port 290 nsew signal input
rlabel metal2 s 259868 -480 259980 240 8 la_oenb[53]
port 291 nsew signal input
rlabel metal2 s 262724 -480 262836 240 8 la_oenb[54]
port 292 nsew signal input
rlabel metal2 s 265580 -480 265692 240 8 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 268436 -480 268548 240 8 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 271292 -480 271404 240 8 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 274148 -480 274260 240 8 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 277004 -480 277116 240 8 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 122780 -480 122892 240 8 la_oenb[5]
port 298 nsew signal input
rlabel metal2 s 279860 -480 279972 240 8 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 282716 -480 282828 240 8 la_oenb[61]
port 300 nsew signal input
rlabel metal2 s 285572 -480 285684 240 8 la_oenb[62]
port 301 nsew signal input
rlabel metal2 s 288428 -480 288540 240 8 la_oenb[63]
port 302 nsew signal input
rlabel metal2 s 125636 -480 125748 240 8 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 128492 -480 128604 240 8 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 131348 -480 131460 240 8 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 134204 -480 134316 240 8 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 289380 -480 289492 240 8 user_clock2
port 307 nsew signal input
rlabel metal2 s 290332 -480 290444 240 8 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 291284 -480 291396 240 8 user_irq[1]
port 309 nsew signal output
rlabel metal2 s 292236 -480 292348 240 8 user_irq[2]
port 310 nsew signal output
rlabel metal4 s -478 -342 -168 298654 4 vdd
port 311 nsew power bidirectional
rlabel metal5 s -478 -342 298510 -32 8 vdd
port 311 nsew power bidirectional
rlabel metal5 s -478 298344 298510 298654 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 298200 -342 298510 298654 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 2709 -822 3019 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 18069 -822 18379 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 33429 -822 33739 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 48789 -822 49099 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 64149 -822 64459 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 79509 -822 79819 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 94869 -822 95179 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 110229 -822 110539 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 125589 -822 125899 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 140949 -822 141259 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 156309 -822 156619 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 171669 -822 171979 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 187029 -822 187339 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 202389 -822 202699 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 217749 -822 218059 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 233109 -822 233419 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 248469 -822 248779 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 263829 -822 264139 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 279189 -822 279499 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 294549 -822 294859 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 1913 298990 2223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 10913 298990 11223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 19913 298990 20223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 28913 298990 29223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 37913 298990 38223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 46913 298990 47223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 55913 298990 56223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 64913 298990 65223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 73913 298990 74223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 82913 298990 83223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 91913 298990 92223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 100913 298990 101223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 109913 298990 110223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 118913 298990 119223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 127913 298990 128223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 136913 298990 137223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 145913 298990 146223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 154913 298990 155223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 163913 298990 164223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 172913 298990 173223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 181913 298990 182223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 190913 298990 191223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 199913 298990 200223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 208913 298990 209223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 217913 298990 218223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 226913 298990 227223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 235913 298990 236223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 244913 298990 245223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 253913 298990 254223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 262913 298990 263223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 271913 298990 272223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 280913 298990 281223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 289913 298990 290223 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s -958 -822 -648 299134 4 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 -822 298990 -512 8 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 298824 298990 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 298680 -822 298990 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 4569 -822 4879 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 19929 -822 20239 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 35289 -822 35599 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 50649 -822 50959 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 66009 -822 66319 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 81369 -822 81679 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 96729 -822 97039 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 112089 -822 112399 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 127449 -822 127759 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 142809 -822 143119 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 158169 -822 158479 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 173529 -822 173839 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 188889 -822 189199 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 204249 -822 204559 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 219609 -822 219919 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 234969 -822 235279 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 250329 -822 250639 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 265689 -822 265999 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 281049 -822 281359 109205 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 281049 112587 281359 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 296409 -822 296719 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 4913 298990 5223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 13913 298990 14223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 22913 298990 23223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 31913 298990 32223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 40913 298990 41223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 49913 298990 50223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 58913 298990 59223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 67913 298990 68223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 76913 298990 77223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 85913 298990 86223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 94913 298990 95223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 103913 298990 104223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 112913 298990 113223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 121913 298990 122223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 130913 298990 131223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 139913 298990 140223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 148913 298990 149223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 157913 298990 158223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 166913 298990 167223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 175913 298990 176223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 184913 298990 185223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 193913 298990 194223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 202913 298990 203223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 211913 298990 212223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 220913 298990 221223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 229913 298990 230223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 238913 298990 239223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 247913 298990 248223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 256913 298990 257223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 265913 298990 266223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 274913 298990 275223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 283913 298990 284223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 292913 298990 293223 6 vss
port 312 nsew ground bidirectional
rlabel metal2 s 5684 -480 5796 240 8 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 6636 -480 6748 240 8 wb_rst_i
port 314 nsew signal input
rlabel metal2 s 7588 -480 7700 240 8 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 11396 -480 11508 240 8 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 43764 -480 43876 240 8 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal2 s 46620 -480 46732 240 8 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 49476 -480 49588 240 8 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 52332 -480 52444 240 8 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal2 s 55188 -480 55300 240 8 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal2 s 58044 -480 58156 240 8 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 60900 -480 61012 240 8 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal2 s 63756 -480 63868 240 8 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal2 s 66612 -480 66724 240 8 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 69468 -480 69580 240 8 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal2 s 15204 -480 15316 240 8 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 72324 -480 72436 240 8 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 75180 -480 75292 240 8 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 78036 -480 78148 240 8 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal2 s 80892 -480 81004 240 8 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 83748 -480 83860 240 8 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal2 s 86604 -480 86716 240 8 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 89460 -480 89572 240 8 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 92316 -480 92428 240 8 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal2 s 95172 -480 95284 240 8 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal2 s 98028 -480 98140 240 8 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 19012 -480 19124 240 8 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal2 s 100884 -480 100996 240 8 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal2 s 103740 -480 103852 240 8 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 22820 -480 22932 240 8 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 26628 -480 26740 240 8 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 29484 -480 29596 240 8 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal2 s 32340 -480 32452 240 8 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 35196 -480 35308 240 8 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 38052 -480 38164 240 8 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal2 s 40908 -480 41020 240 8 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 8540 -480 8652 240 8 wbs_cyc_i
port 348 nsew signal input
rlabel metal2 s 12348 -480 12460 240 8 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal2 s 44716 -480 44828 240 8 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 47572 -480 47684 240 8 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal2 s 50428 -480 50540 240 8 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 53284 -480 53396 240 8 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal2 s 56140 -480 56252 240 8 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal2 s 58996 -480 59108 240 8 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 61852 -480 61964 240 8 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 64708 -480 64820 240 8 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 67564 -480 67676 240 8 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 70420 -480 70532 240 8 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 16156 -480 16268 240 8 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal2 s 73276 -480 73388 240 8 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 76132 -480 76244 240 8 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal2 s 78988 -480 79100 240 8 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal2 s 81844 -480 81956 240 8 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal2 s 84700 -480 84812 240 8 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 87556 -480 87668 240 8 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 90412 -480 90524 240 8 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 93268 -480 93380 240 8 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 96124 -480 96236 240 8 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal2 s 98980 -480 99092 240 8 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 19964 -480 20076 240 8 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal2 s 101836 -480 101948 240 8 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal2 s 104692 -480 104804 240 8 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 23772 -480 23884 240 8 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 27580 -480 27692 240 8 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 30436 -480 30548 240 8 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal2 s 33292 -480 33404 240 8 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 36148 -480 36260 240 8 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal2 s 39004 -480 39116 240 8 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 41860 -480 41972 240 8 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal2 s 13300 -480 13412 240 8 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal2 s 45668 -480 45780 240 8 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 48524 -480 48636 240 8 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal2 s 51380 -480 51492 240 8 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 54236 -480 54348 240 8 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 57092 -480 57204 240 8 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 59948 -480 60060 240 8 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal2 s 62804 -480 62916 240 8 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal2 s 65660 -480 65772 240 8 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 68516 -480 68628 240 8 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 71372 -480 71484 240 8 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 17108 -480 17220 240 8 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal2 s 74228 -480 74340 240 8 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 77084 -480 77196 240 8 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 79940 -480 80052 240 8 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal2 s 82796 -480 82908 240 8 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 85652 -480 85764 240 8 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 88508 -480 88620 240 8 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 91364 -480 91476 240 8 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 94220 -480 94332 240 8 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 97076 -480 97188 240 8 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 99932 -480 100044 240 8 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal2 s 20916 -480 21028 240 8 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal2 s 102788 -480 102900 240 8 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal2 s 105644 -480 105756 240 8 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 24724 -480 24836 240 8 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 28532 -480 28644 240 8 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal2 s 31388 -480 31500 240 8 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal2 s 34244 -480 34356 240 8 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 37100 -480 37212 240 8 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 39956 -480 40068 240 8 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 42812 -480 42924 240 8 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 14252 -480 14364 240 8 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 18060 -480 18172 240 8 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 21868 -480 21980 240 8 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal2 s 25676 -480 25788 240 8 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal2 s 9492 -480 9604 240 8 wbs_stb_i
port 417 nsew signal input
rlabel metal2 s 10444 -480 10556 240 8 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 298020 298020
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17260670
string GDS_FILE /mnt/c/Users/aidan/caravel_user_project/openlane/user_project_wrapper/runs/23_12_10_16_56/results/signoff/user_project_wrapper.magic.gds
string GDS_START 15160638
<< end >>

