magic
tech gf180mcuD
magscale 1 5
timestamp 1702242473
<< obsm1 >>
rect 672 1538 279328 174078
<< metal2 >>
rect 139888 0 139944 400
<< obsm2 >>
rect 854 430 279202 174067
rect 854 400 139858 430
rect 139974 400 279202 430
<< metal3 >>
rect 279600 169456 280000 169512
rect 279600 156912 280000 156968
rect 279600 144368 280000 144424
rect 279600 131824 280000 131880
rect 279600 119280 280000 119336
rect 279600 106736 280000 106792
rect 279600 94192 280000 94248
rect 0 87920 400 87976
rect 279600 81648 280000 81704
rect 279600 69104 280000 69160
rect 279600 56560 280000 56616
rect 279600 44016 280000 44072
rect 279600 31472 280000 31528
rect 279600 18928 280000 18984
rect 279600 6384 280000 6440
<< obsm3 >>
rect 400 169542 279600 174062
rect 400 169426 279570 169542
rect 400 156998 279600 169426
rect 400 156882 279570 156998
rect 400 144454 279600 156882
rect 400 144338 279570 144454
rect 400 131910 279600 144338
rect 400 131794 279570 131910
rect 400 119366 279600 131794
rect 400 119250 279570 119366
rect 400 106822 279600 119250
rect 400 106706 279570 106822
rect 400 94278 279600 106706
rect 400 94162 279570 94278
rect 400 88006 279600 94162
rect 430 87890 279600 88006
rect 400 81734 279600 87890
rect 400 81618 279570 81734
rect 400 69190 279600 81618
rect 400 69074 279570 69190
rect 400 56646 279600 69074
rect 400 56530 279570 56646
rect 400 44102 279600 56530
rect 400 43986 279570 44102
rect 400 31558 279600 43986
rect 400 31442 279570 31558
rect 400 19014 279600 31442
rect 400 18898 279570 19014
rect 400 6470 279600 18898
rect 400 6354 279570 6470
rect 400 1554 279600 6354
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< obsm4 >>
rect 279062 108761 279090 110031
<< labels >>
rlabel metal3 s 279600 6384 280000 6440 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 279600 44016 280000 44072 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 279600 81648 280000 81704 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 279600 119280 280000 119336 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 279600 131824 280000 131880 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 279600 144368 280000 144424 6 io_in[5]
port 6 nsew signal input
rlabel metal3 s 279600 156912 280000 156968 6 io_in[6]
port 7 nsew signal input
rlabel metal3 s 279600 169456 280000 169512 6 io_in[7]
port 8 nsew signal input
rlabel metal3 s 0 87920 400 87976 6 io_in[8]
port 9 nsew signal input
rlabel metal3 s 279600 31472 280000 31528 6 io_oeb[0]
port 10 nsew signal output
rlabel metal3 s 279600 69104 280000 69160 6 io_oeb[1]
port 11 nsew signal output
rlabel metal3 s 279600 106736 280000 106792 6 io_oeb[2]
port 12 nsew signal output
rlabel metal3 s 279600 18928 280000 18984 6 io_out[0]
port 13 nsew signal output
rlabel metal3 s 279600 56560 280000 56616 6 io_out[1]
port 14 nsew signal output
rlabel metal3 s 279600 94192 280000 94248 6 io_out[2]
port 15 nsew signal output
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 17 nsew ground bidirectional
rlabel metal2 s 139888 0 139944 400 6 wb_clk_i
port 18 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15160584
string GDS_FILE /mnt/c/Users/aidan/caravel_user_project/openlane/user_proj_example/runs/23_12_10_15_47/results/signoff/user_proj_example.magic.gds
string GDS_START 202120
<< end >>

